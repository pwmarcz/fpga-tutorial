module counter(input wire       clk,
               input wire       en,
               input wire       rst,
               output reg [3:0] count);
  // TODO
endmodule
