module traffic(input wire  clk,
               input wire  go,
               output wire red,
               output wire yellow,
               output wire green);
  // TODO
endmodule
