module serial(input wire clk,
              input wire in,
              input wire [7:0] data,
              output wire ready,
              output wire out);
  // TODO
endmodule
